`include "GUVM_test.sv"
`include"add_test.sv"
`include"bie_test.sv"
`include"child_test.sv"