`include "GUVM_test.sv"
`include"add_test.sv"
`include"bie_test.sv"