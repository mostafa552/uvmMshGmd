`include "add.svh"
`include "test.svh"
`include "jal.svh"
`include "load.svh"
`include "store.svh"
`include "nop.svh"
`include "addcc.svh"
`include "addx.svh"
`include "bie.svh"
`include "ba.svh"